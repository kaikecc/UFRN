library verilog;
use verilog.vl_types.all;
entity mux8x1_vlg_check_tst is
    port(
        M8              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux8x1_vlg_check_tst;
