library verilog;
use verilog.vl_types.all;
entity MUX_Display_vlg_check_tst is
    port(
        MD              : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end MUX_Display_vlg_check_tst;
