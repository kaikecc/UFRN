library verilog;
use verilog.vl_types.all;
entity MUX_comp1_vlg_vec_tst is
end MUX_comp1_vlg_vec_tst;
