library verilog;
use verilog.vl_types.all;
entity mux8x1_vlg_vec_tst is
end mux8x1_vlg_vec_tst;
