library verilog;
use verilog.vl_types.all;
entity REGS_GRV_vlg_vec_tst is
end REGS_GRV_vlg_vec_tst;
