ENTITY BITCOMPARADOR IS
	PORT( A,B,AM,BM,ABIG : IN BIT;
	AB,BA,IG : OUT BIT);
END BITCOMPARADOR;

ARCHITECTURE CKT OF BITCOMPARADOR IS

BEGIN
  AB<=(A AND NOT B AND ABIG) OR (AM);
  BA<=(B AND NOT A AND ABIG) OR (BM);
  IG<=ABIG AND (A XNOR B);
END CKT ;





