library verilog;
use verilog.vl_types.all;
entity Comparador_vlg_vec_tst is
end Comparador_vlg_vec_tst;
