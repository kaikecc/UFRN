library verilog;
use verilog.vl_types.all;
entity MUX2_comp1_vlg_vec_tst is
end MUX2_comp1_vlg_vec_tst;
