library verilog;
use verilog.vl_types.all;
entity reg8bit_vlg_vec_tst is
end reg8bit_vlg_vec_tst;
