library verilog;
use verilog.vl_types.all;
entity MUX1_comp1_vlg_vec_tst is
end MUX1_comp1_vlg_vec_tst;
