library verilog;
use verilog.vl_types.all;
entity mde_vlg_vec_tst is
end mde_vlg_vec_tst;
