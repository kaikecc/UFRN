library verilog;
use verilog.vl_types.all;
entity MUX_SUM_vlg_vec_tst is
end MUX_SUM_vlg_vec_tst;
