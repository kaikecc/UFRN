library verilog;
use verilog.vl_types.all;
entity somador8bit_vlg_vec_tst is
end somador8bit_vlg_vec_tst;
