library verilog;
use verilog.vl_types.all;
entity multiplicador4bit_vlg_vec_tst is
end multiplicador4bit_vlg_vec_tst;
