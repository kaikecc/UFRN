library verilog;
use verilog.vl_types.all;
entity subtrator8bit_vlg_vec_tst is
end subtrator8bit_vlg_vec_tst;
