library verilog;
use verilog.vl_types.all;
entity comparador4bit_vlg_vec_tst is
end comparador4bit_vlg_vec_tst;
