library verilog;
use verilog.vl_types.all;
entity contador8bit_vlg_vec_tst is
end contador8bit_vlg_vec_tst;
