library verilog;
use verilog.vl_types.all;
entity comparador8bit_vlg_vec_tst is
end comparador8bit_vlg_vec_tst;
