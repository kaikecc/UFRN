library verilog;
use verilog.vl_types.all;
entity mde is
    port(
        ck              : in     vl_logic;
        b_on            : in     vl_logic;
        b_next          : in     vl_logic;
        b_back          : in     vl_logic;
        play            : in     vl_logic;
        cont_local_10   : in     vl_logic;
        cont_on_5       : in     vl_logic;
        it_comparador   : in     vl_logic;
        grt_comparador  : in     vl_logic;
        eq_comparador   : in     vl_logic;
        nova_msg        : in     vl_logic;
        F_led           : out    vl_logic;
        M_led           : out    vl_logic;
        P_led           : out    vl_logic;
        O_led           : out    vl_logic;
        R_led           : out    vl_logic;
        ld_display_val  : out    vl_logic;
        r_w             : out    vl_logic;
        en              : out    vl_logic;
        DISPLAY_EN      : out    vl_logic;
        sub_display     : out    vl_logic;
        erase_MEM       : out    vl_logic;
        sum_Display     : out    vl_logic;
        clr_addr        : out    vl_logic;
        setUni          : out    vl_logic;
        sl_comp1        : out    vl_logic;
        sl1_comp1       : out    vl_logic;
        sl2_comp1       : out    vl_logic;
        s_comp1         : out    vl_logic;
        s1_comp1        : out    vl_logic;
        s2_comp1        : out    vl_logic;
        clr_Cont_local  : out    vl_logic;
        clr_CT_ON       : out    vl_logic;
        clr_CT_Msg      : out    vl_logic;
        clr_CT_INAT     : out    vl_logic;
        en_CT_INAT      : out    vl_logic;
        en_Cont_local   : out    vl_logic;
        en_CT_Msg       : out    vl_logic;
        en_CT_ON        : out    vl_logic;
        ld_REGS_REP_SQ  : out    vl_logic;
        ld_REGS_REP_S   : out    vl_logic;
        ld_REGS_GRV     : out    vl_logic;
        Flag_rep_s      : out    vl_logic;
        Flag_rep_sq     : out    vl_logic;
        clr_REGS_REP    : out    vl_logic
    );
end mde;
