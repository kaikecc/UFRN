library verilog;
use verilog.vl_types.all;
entity multiplicador8bit_vlg_vec_tst is
end multiplicador8bit_vlg_vec_tst;
