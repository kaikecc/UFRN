library verilog;
use verilog.vl_types.all;
entity CT_Msg_vlg_vec_tst is
end CT_Msg_vlg_vec_tst;
