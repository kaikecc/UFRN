library verilog;
use verilog.vl_types.all;
entity MUX_Display_vlg_vec_tst is
end MUX_Display_vlg_vec_tst;
